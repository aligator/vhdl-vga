../vga_sync_gen/vga_sync_gen.vhdl